--vhdl1
